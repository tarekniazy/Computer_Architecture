
Library ieee;
use ieee.std_Logic_1164.all;

ENTITY Control is 
  PORT ( Opcode : IN std_logic_vector (4 DOWNTO 0);
         clk,Interrupt :  IN std_logic;
         Reset :  IN std_logic;
         Signals : OUT std_logic_vector (0 TO 38);
         Zf,Cf,Nf: OUT std_logic;
           ldm_in :OUT std_logic);  
  END Control;
  
  ARCHITECTURE a_Control OF Control
  IS 
    type Op_Array is array (0 to 27) of std_logic_vector (4 DOWNTO 0);    
    type Signalm_Array is array (0 to 4) of std_logic_vector (0 TO 38);
    type Signalj_Array is array (0 to 6) of std_logic_vector (0 TO 38);
    type Signal_Array is array (0 to 7) of std_logic_vector (0 TO 38);
    signal Opcode_s : Op_Array := ("00000","00001","00010","00011","00100","00101","00110","00111","01000","01001","01010","01011","01100","01101","01110","01111","10000","10001","10010","10011","10100","10101","10110","10111","11000","11001","11010","11011");
    signal Signals_one : Signal_Array  := ("000000000000000000000000000000001111100","000001100000000001010000011000001111100","000001100000000001011000011000001111100","000011100000010000111100011000001111100","000011100000010000000100011000001111100","000011100000010000011100011000001111100","000011100000000000000000001100001111100","000011100000001000110100001000001111101");   
 --signal Signals_one : Signal_Array  := ("0000000000000000000000000000000011111","0000011000000000010100000110000011111","0000011000000000010110000110000011111","0000111000000100001111000110000011111","0000111000000100000001000110000011111","0000111000000100000111000110000011111","0000111000000000000000000011000011111","0000111000000010000001000010000011111");
      signal Signals_two : Signal_Array  := ("000001100000000100000110001000001111100","001101101000010000001100011000001111100","000001110000010000001100011000001111100","000101101000010000010100011000001111100","000101101000010000100100011000001111100","000101101000010000101100011000001111100","000011100100010001001100011000001111100","000011100100010001000100011000001111100");
 --signal Signals_two : Signal_Array  := ("0000011000000001000001100010000011111","0001011000000001000001000110000011111","0000011100000100000011000110000011111","0001011010000100000101000110000011111","0001011010000100001001000110000011111","0001011010000100001011000110000011111","0000111001000100010011000110000011111","0000111001000100010001000110000011111");
    signal Signals_mem : Signalm_Array := ("000001100001000000000000101011101111100","000011100000000010000101001000101111100","000011110000010000110100001000001111100","000011100010000000110101001000001111100","000001100011000000110000101000001111100");
    signal Signals_jmp : Signalj_Array := ("100000000000000000000000001000001110000","100000100000000000000000001000001110000","100001000000000000000000001000001110000","100000000000000000000000001000011110000","100000000000000000000000111011111111000","100000000000000010000001011001101111110","100000000000000010000001011001111111100");
    BEGIN
  
  process (Opcode,Reset,Interrupt,clk)
    begin

 IF Opcode = "10101" THEN
      Zf <= '1';
      Cf <= '0';
      Nf <= '0';

  ELSIF Opcode = "10110" THEN
      Zf <= '0';
      Cf <= '0';
      Nf <= '1';

  ELSIF Opcode = "10111" THEN
      Zf <= '0';
      Cf <= '1';
      Nf <= '0';
  ELSE 
     Zf <= '0';
     Cf <= '0';
     Nf <= '0';
  END IF;
--if rising_edge(clk) then
  IF (Reset = '0') and (Interrupt ='0') THEN
    For i in 0 to 7 Loop
      IF Opcode = Opcode_s(i) THEN
        Signals <= Signals_one(i);     
      END IF;    
    end loop;
    For i in 8 to 15 Loop
      IF Opcode = Opcode_s(i) THEN
        Signals <= Signals_two(i-8);     
      END IF;    
    end loop;
    For i in 16 to 20 Loop
      IF Opcode = Opcode_s(i) THEN
        Signals <= Signals_mem(i-16);     
      END IF;    
    end loop;
    For i in 21 to 27 Loop
      IF Opcode = Opcode_s(i) THEN
        Signals <= Signals_jmp(i-21);     
      END IF;    
    end loop;
  END IF;
 --end if;
if Opcode = "10010" THEN

ldm_in<='1';

else 

ldm_in<='0';


end if;

end process;
  END a_Control;